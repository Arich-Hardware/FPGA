------------------------------------------------------------------------
-- trig_tdc.vhd
--
-- trigger input TDC
------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.tdc_types.all;

entity trigger_tdc_with_fifo is

  port (
    clk         : in  std_logic_vector(3 downto 0);  -- 4 phase clock
    rst         : in  std_logic;                     -- active high asynch
    trigger     : in  std_logic;                     -- rising edge
    empty, full : out std_logic;
    output      : out trigger_tdc_hit;               -- hit (time, phase, evn)
    rd_ena      : in  std_logic);

end entity trigger_tdc_with_fifo;

architecture synth of trigger_tdc_with_fifo is

  component trigger_tdc is
    port (
      clk          : in  std_logic_vector(3 downto 0);
      rst          : in  std_logic;
      trigger      : in  std_logic;
      output       : out trigger_tdc_hit;
      output_valid : out std_logic);
  end component trigger_tdc;

  component web_fifo is
    generic (
      RAM_WIDTH : natural;
      RAM_DEPTH : natural);
    port (
      clk        : in  std_logic;
      rst        : in  std_logic;
      wr_en      : in  std_logic;
      wr_data    : in  std_logic_vector(RAM_WIDTH - 1 downto 0);
      rd_en      : in  std_logic;
      rd_valid   : out std_logic;
      rd_data    : out std_logic_vector(RAM_WIDTH - 1 downto 0);
      empty      : out std_logic;
      empty_next : out std_logic;
      full       : out std_logic;
      full_next  : out std_logic;
      fill_count : out integer range RAM_DEPTH - 1 downto 0);
  end component web_fifo;

  signal trigger_data : trigger_tdc_hit;
  signal trigger_data_v : std_logic_vector( len(trigger_data)-1 downto 0);
  signal trigger_valid : std_logic;

  signal output_data : trigger_tdc_hit;
  signal output_data_v : std_logic_vector( len(output_data)-1 downto 0);

begin  -- architecture synth

  trigger_tdc_1: entity work.trigger_tdc
    port map (
      clk          => clk,
      rst          => rst,
      trigger      => trigger,
      output       => trigger_data,
      output_valid => trigger_valid);

  web_fifo_1: entity work.web_fifo
    generic map (
      RAM_WIDTH => len( output_data_v),
      RAM_DEPTH => 16)
    port map (
      clk        => clk(0),
      rst        => rst,
      wr_en      => trigger_valid,
      wr_data    => trigger_data_v,
      rd_en      => rd_ena,
      rd_valid   => open,
      rd_data    => output_data_v,
      empty      => empty,
      empty_next => open,
      full       => full,
      full_next  => open,
      fill_count => open);

  trigger_data_v <= vectorify( trigger_data, trigger_data_v);
  output_data <= structify( output_data_v, output_data);

  output <= output_data;

end architecture synth;
